-- 32-bit Adder
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity cacheC is
    port (instruction : in bit_vector(31 downto 0);
    tag : in bit_vector(9 downto 0));
end cacheC;

architecture behave of cacheC is
begin  -- behave
    
    

end behave;

